package MIPSCPU_constants is
--set to 31 instead of 32 to accomodate 0th bit
constant register_size : integer := 31;
end MIPSCPU_constants;